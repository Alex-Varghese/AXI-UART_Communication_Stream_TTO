QuestaSim vlog 10.6c Compiler 2017.07 Jul 25 2017
Start time: 15:42:04 on Nov 04,2025
vlog -sv "+acc" "+cover" "+fcover" -l package.sv top.sv 
-- Compiling module uart_rec
-- Compiling module uart_tx
-- Compiling module sync_fifo
-- Compiling module axis_fifo_uart_tx
-- Compiling module axis_master_inp
-- Compiling module top_axis_uart
-- Compiling interface intf
-- Compiling module assertions
-- Compiling package top_sv_unit
-- Importing package mtiUvm.uvm_pkg (uvm-1.1d Built-in)
-- Importing package pkg
-- Compiling module top

Top level modules:
	assertions
	top
End time: 15:42:05 on Nov 04,2025, Elapsed time: 0:00:01
Errors: 0, Warnings: 0
